module sine_rom( input  logic                clk,
                 input  logic unsigned [7:0] addr,
                 output logic unsigned [7:0] val );

    always_ff @(posedge clk)
        case(addr)
                0 : val <= 127;
                1 : val <= 127;
                2 : val <= 128;
                3 : val <= 128;
                4 : val <= 129;
                5 : val <= 129;
                6 : val <= 129;
                7 : val <= 130;
                8 : val <= 130;
                9 : val <= 131;
                10 : val <= 131;
                11 : val <= 131;
                12 : val <= 132;
                13 : val <= 132;
                14 : val <= 132;
                15 : val <= 133;
                16 : val <= 133;
                17 : val <= 134;
                18 : val <= 134;
                19 : val <= 134;
                20 : val <= 135;
                21 : val <= 135;
                22 : val <= 136;
                23 : val <= 136;
                24 : val <= 136;
                25 : val <= 137;
                26 : val <= 137;
                27 : val <= 138;
                28 : val <= 138;
                29 : val <= 138;
                30 : val <= 139;
                31 : val <= 139;
                32 : val <= 139;
                33 : val <= 140;
                34 : val <= 140;
                35 : val <= 141;
                36 : val <= 141;
                37 : val <= 141;
                38 : val <= 142;
                39 : val <= 142;
                40 : val <= 143;
                41 : val <= 143;
                42 : val <= 143;
                43 : val <= 144;
                44 : val <= 144;
                45 : val <= 145;
                46 : val <= 145;
                47 : val <= 145;
                48 : val <= 146;
                49 : val <= 146;
                50 : val <= 146;
                51 : val <= 147;
                52 : val <= 147;
                53 : val <= 148;
                54 : val <= 148;
                55 : val <= 148;
                56 : val <= 149;
                57 : val <= 149;
                58 : val <= 150;
                59 : val <= 150;
                60 : val <= 150;
                61 : val <= 151;
                62 : val <= 151;
                63 : val <= 151;
                64 : val <= 152;
                65 : val <= 152;
                66 : val <= 153;
                67 : val <= 153;
                68 : val <= 153;
                69 : val <= 154;
                70 : val <= 154;
                71 : val <= 155;
                72 : val <= 155;
                73 : val <= 155;
                74 : val <= 156;
                75 : val <= 156;
                76 : val <= 156;
                77 : val <= 157;
                78 : val <= 157;
                79 : val <= 158;
                80 : val <= 158;
                81 : val <= 158;
                82 : val <= 159;
                83 : val <= 159;
                84 : val <= 159;
                85 : val <= 160;
                86 : val <= 160;
                87 : val <= 161;
                88 : val <= 161;
                89 : val <= 161;
                90 : val <= 162;
                91 : val <= 162;
                92 : val <= 163;
                93 : val <= 163;
                94 : val <= 163;
                95 : val <= 164;
                96 : val <= 164;
                97 : val <= 164;
                98 : val <= 165;
                99 : val <= 165;
                100 : val <= 166;
                101 : val <= 166;
                102 : val <= 166;
                103 : val <= 167;
                104 : val <= 167;
                105 : val <= 167;
                106 : val <= 168;
                107 : val <= 168;
                108 : val <= 168;
                109 : val <= 169;
                110 : val <= 169;
                111 : val <= 170;
                112 : val <= 170;
                113 : val <= 170;
                114 : val <= 171;
                115 : val <= 171;
                116 : val <= 171;
                117 : val <= 172;
                118 : val <= 172;
                119 : val <= 173;
                120 : val <= 173;
                121 : val <= 173;
                122 : val <= 174;
                123 : val <= 174;
                124 : val <= 174;
                125 : val <= 175;
                126 : val <= 175;
                127 : val <= 175;
                128 : val <= 176;
                129 : val <= 176;
                130 : val <= 177;
                131 : val <= 177;
                132 : val <= 177;
                133 : val <= 178;
                134 : val <= 178;
                135 : val <= 178;
                136 : val <= 179;
                137 : val <= 179;
                138 : val <= 179;
                139 : val <= 180;
                140 : val <= 180;
                141 : val <= 180;
                142 : val <= 181;
                143 : val <= 181;
                144 : val <= 182;
                145 : val <= 182;
                146 : val <= 182;
                147 : val <= 183;
                148 : val <= 183;
                149 : val <= 183;
                150 : val <= 184;
                151 : val <= 184;
                152 : val <= 184;
                153 : val <= 185;
                154 : val <= 185;
                155 : val <= 185;
                156 : val <= 186;
                157 : val <= 186;
                158 : val <= 186;
                159 : val <= 187;
                160 : val <= 187;
                161 : val <= 187;
                162 : val <= 188;
                163 : val <= 188;
                164 : val <= 188;
                165 : val <= 189;
                166 : val <= 189;
                167 : val <= 190;
                168 : val <= 190;
                169 : val <= 190;
                170 : val <= 191;
                171 : val <= 191;
                172 : val <= 191;
                173 : val <= 192;
                174 : val <= 192;
                175 : val <= 192;
                176 : val <= 193;
                177 : val <= 193;
                178 : val <= 193;
                179 : val <= 194;
                180 : val <= 194;
                181 : val <= 194;
                182 : val <= 195;
                183 : val <= 195;
                184 : val <= 195;
                185 : val <= 196;
                186 : val <= 196;
                187 : val <= 196;
                188 : val <= 197;
                189 : val <= 197;
                190 : val <= 197;
                191 : val <= 198;
                192 : val <= 198;
                193 : val <= 198;
                194 : val <= 198;
                195 : val <= 199;
                196 : val <= 199;
                197 : val <= 199;
                198 : val <= 200;
                199 : val <= 200;
                200 : val <= 200;
                201 : val <= 201;
                202 : val <= 201;
                203 : val <= 201;
                204 : val <= 202;
                205 : val <= 202;
                206 : val <= 202;
                207 : val <= 203;
                208 : val <= 203;
                209 : val <= 203;
                210 : val <= 204;
                211 : val <= 204;
                212 : val <= 204;
                213 : val <= 205;
                214 : val <= 205;
                215 : val <= 205;
                216 : val <= 205;
                217 : val <= 206;
                218 : val <= 206;
                219 : val <= 206;
                220 : val <= 207;
                221 : val <= 207;
                222 : val <= 207;
                223 : val <= 208;
                224 : val <= 208;
                225 : val <= 208;
                226 : val <= 208;
                227 : val <= 209;
                228 : val <= 209;
                229 : val <= 209;
                230 : val <= 210;
                231 : val <= 210;
                232 : val <= 210;
                233 : val <= 211;
                234 : val <= 211;
                235 : val <= 211;
                236 : val <= 211;
                237 : val <= 212;
                238 : val <= 212;
                239 : val <= 212;
                240 : val <= 213;
                241 : val <= 213;
                242 : val <= 213;
                243 : val <= 213;
                244 : val <= 214;
                245 : val <= 214;
                246 : val <= 214;
                247 : val <= 215;
                248 : val <= 215;
                249 : val <= 215;
                250 : val <= 215;
                251 : val <= 216;
                252 : val <= 216;
                253 : val <= 216;
                254 : val <= 217;
                255 : val <= 217;
                256 : val <= 217;
                257 : val <= 217;
                258 : val <= 218;
                259 : val <= 218;
                260 : val <= 218;
                261 : val <= 219;
                262 : val <= 219;
                263 : val <= 219;
                264 : val <= 219;
                265 : val <= 220;
                266 : val <= 220;
                267 : val <= 220;
                268 : val <= 220;
                269 : val <= 221;
                270 : val <= 221;
                271 : val <= 221;
                272 : val <= 221;
                273 : val <= 222;
                274 : val <= 222;
                275 : val <= 222;
                276 : val <= 223;
                277 : val <= 223;
                278 : val <= 223;
                279 : val <= 223;
                280 : val <= 224;
                281 : val <= 224;
                282 : val <= 224;
                283 : val <= 224;
                284 : val <= 225;
                285 : val <= 225;
                286 : val <= 225;
                287 : val <= 225;
                288 : val <= 226;
                289 : val <= 226;
                290 : val <= 226;
                291 : val <= 226;
                292 : val <= 227;
                293 : val <= 227;
                294 : val <= 227;
                295 : val <= 227;
                296 : val <= 228;
                297 : val <= 228;
                298 : val <= 228;
                299 : val <= 228;
                300 : val <= 228;
                301 : val <= 229;
                302 : val <= 229;
                303 : val <= 229;
                304 : val <= 229;
                305 : val <= 230;
                306 : val <= 230;
                307 : val <= 230;
                308 : val <= 230;
                309 : val <= 231;
                310 : val <= 231;
                311 : val <= 231;
                312 : val <= 231;
                313 : val <= 231;
                314 : val <= 232;
                315 : val <= 232;
                316 : val <= 232;
                317 : val <= 232;
                318 : val <= 233;
                319 : val <= 233;
                320 : val <= 233;
                321 : val <= 233;
                322 : val <= 233;
                323 : val <= 234;
                324 : val <= 234;
                325 : val <= 234;
                326 : val <= 234;
                327 : val <= 235;
                328 : val <= 235;
                329 : val <= 235;
                330 : val <= 235;
                331 : val <= 235;
                332 : val <= 236;
                333 : val <= 236;
                334 : val <= 236;
                335 : val <= 236;
                336 : val <= 236;
                337 : val <= 237;
                338 : val <= 237;
                339 : val <= 237;
                340 : val <= 237;
                341 : val <= 237;
                342 : val <= 238;
                343 : val <= 238;
                344 : val <= 238;
                345 : val <= 238;
                346 : val <= 238;
                347 : val <= 239;
                348 : val <= 239;
                349 : val <= 239;
                350 : val <= 239;
                351 : val <= 239;
                352 : val <= 239;
                353 : val <= 240;
                354 : val <= 240;
                355 : val <= 240;
                356 : val <= 240;
                357 : val <= 240;
                358 : val <= 241;
                359 : val <= 241;
                360 : val <= 241;
                361 : val <= 241;
                362 : val <= 241;
                363 : val <= 241;
                364 : val <= 242;
                365 : val <= 242;
                366 : val <= 242;
                367 : val <= 242;
                368 : val <= 242;
                369 : val <= 242;
                370 : val <= 243;
                371 : val <= 243;
                372 : val <= 243;
                373 : val <= 243;
                374 : val <= 243;
                375 : val <= 243;
                376 : val <= 244;
                377 : val <= 244;
                378 : val <= 244;
                379 : val <= 244;
                380 : val <= 244;
                381 : val <= 244;
                382 : val <= 244;
                383 : val <= 245;
                384 : val <= 245;
                385 : val <= 245;
                386 : val <= 245;
                387 : val <= 245;
                388 : val <= 245;
                389 : val <= 246;
                390 : val <= 246;
                391 : val <= 246;
                392 : val <= 246;
                393 : val <= 246;
                394 : val <= 246;
                395 : val <= 246;
                396 : val <= 247;
                397 : val <= 247;
                398 : val <= 247;
                399 : val <= 247;
                400 : val <= 247;
                401 : val <= 247;
                402 : val <= 247;
                403 : val <= 247;
                404 : val <= 248;
                405 : val <= 248;
                406 : val <= 248;
                407 : val <= 248;
                408 : val <= 248;
                409 : val <= 248;
                410 : val <= 248;
                411 : val <= 248;
                412 : val <= 249;
                413 : val <= 249;
                414 : val <= 249;
                415 : val <= 249;
                416 : val <= 249;
                417 : val <= 249;
                418 : val <= 249;
                419 : val <= 249;
                420 : val <= 249;
                421 : val <= 250;
                422 : val <= 250;
                423 : val <= 250;
                424 : val <= 250;
                425 : val <= 250;
                426 : val <= 250;
                427 : val <= 250;
                428 : val <= 250;
                429 : val <= 250;
                430 : val <= 250;
                431 : val <= 251;
                432 : val <= 251;
                433 : val <= 251;
                434 : val <= 251;
                435 : val <= 251;
                436 : val <= 251;
                437 : val <= 251;
                438 : val <= 251;
                439 : val <= 251;
                440 : val <= 251;
                441 : val <= 251;
                442 : val <= 252;
                443 : val <= 252;
                444 : val <= 252;
                445 : val <= 252;
                446 : val <= 252;
                447 : val <= 252;
                448 : val <= 252;
                449 : val <= 252;
                450 : val <= 252;
                451 : val <= 252;
                452 : val <= 252;
                453 : val <= 252;
                454 : val <= 252;
                455 : val <= 253;
                456 : val <= 253;
                457 : val <= 253;
                458 : val <= 253;
                459 : val <= 253;
                460 : val <= 253;
                461 : val <= 253;
                462 : val <= 253;
                463 : val <= 253;
                464 : val <= 253;
                465 : val <= 253;
                466 : val <= 253;
                467 : val <= 253;
                468 : val <= 253;
                469 : val <= 253;
                470 : val <= 253;
                471 : val <= 253;
                472 : val <= 254;
                473 : val <= 254;
                474 : val <= 254;
                475 : val <= 254;
                476 : val <= 254;
                477 : val <= 254;
                478 : val <= 254;
                479 : val <= 254;
                480 : val <= 254;
                481 : val <= 254;
                482 : val <= 254;
                483 : val <= 254;
                484 : val <= 254;
                485 : val <= 254;
                486 : val <= 254;
                487 : val <= 254;
                488 : val <= 254;
                489 : val <= 254;
                490 : val <= 254;
                491 : val <= 254;
                492 : val <= 254;
                493 : val <= 254;
                494 : val <= 254;
                495 : val <= 254;
                496 : val <= 254;
                497 : val <= 254;
                498 : val <= 254;
                499 : val <= 254;
                500 : val <= 254;
                501 : val <= 254;
                502 : val <= 254;
                503 : val <= 254;
                504 : val <= 254;
                505 : val <= 254;
                506 : val <= 254;
                507 : val <= 254;
                508 : val <= 254;
                509 : val <= 254;
                510 : val <= 254;
                511 : val <= 254;
                512 : val <= 255;
                513 : val <= 254;
                514 : val <= 254;
                515 : val <= 254;
                516 : val <= 254;
                517 : val <= 254;
                518 : val <= 254;
                519 : val <= 254;
                520 : val <= 254;
                521 : val <= 254;
                522 : val <= 254;
                523 : val <= 254;
                524 : val <= 254;
                525 : val <= 254;
                526 : val <= 254;
                527 : val <= 254;
                528 : val <= 254;
                529 : val <= 254;
                530 : val <= 254;
                531 : val <= 254;
                532 : val <= 254;
                533 : val <= 254;
                534 : val <= 254;
                535 : val <= 254;
                536 : val <= 254;
                537 : val <= 254;
                538 : val <= 254;
                539 : val <= 254;
                540 : val <= 254;
                541 : val <= 254;
                542 : val <= 254;
                543 : val <= 254;
                544 : val <= 254;
                545 : val <= 254;
                546 : val <= 254;
                547 : val <= 254;
                548 : val <= 254;
                549 : val <= 254;
                550 : val <= 254;
                551 : val <= 254;
                552 : val <= 254;
                553 : val <= 253;
                554 : val <= 253;
                555 : val <= 253;
                556 : val <= 253;
                557 : val <= 253;
                558 : val <= 253;
                559 : val <= 253;
                560 : val <= 253;
                561 : val <= 253;
                562 : val <= 253;
                563 : val <= 253;
                564 : val <= 253;
                565 : val <= 253;
                566 : val <= 253;
                567 : val <= 253;
                568 : val <= 253;
                569 : val <= 253;
                570 : val <= 252;
                571 : val <= 252;
                572 : val <= 252;
                573 : val <= 252;
                574 : val <= 252;
                575 : val <= 252;
                576 : val <= 252;
                577 : val <= 252;
                578 : val <= 252;
                579 : val <= 252;
                580 : val <= 252;
                581 : val <= 252;
                582 : val <= 252;
                583 : val <= 251;
                584 : val <= 251;
                585 : val <= 251;
                586 : val <= 251;
                587 : val <= 251;
                588 : val <= 251;
                589 : val <= 251;
                590 : val <= 251;
                591 : val <= 251;
                592 : val <= 251;
                593 : val <= 251;
                594 : val <= 250;
                595 : val <= 250;
                596 : val <= 250;
                597 : val <= 250;
                598 : val <= 250;
                599 : val <= 250;
                600 : val <= 250;
                601 : val <= 250;
                602 : val <= 250;
                603 : val <= 250;
                604 : val <= 249;
                605 : val <= 249;
                606 : val <= 249;
                607 : val <= 249;
                608 : val <= 249;
                609 : val <= 249;
                610 : val <= 249;
                611 : val <= 249;
                612 : val <= 249;
                613 : val <= 248;
                614 : val <= 248;
                615 : val <= 248;
                616 : val <= 248;
                617 : val <= 248;
                618 : val <= 248;
                619 : val <= 248;
                620 : val <= 248;
                621 : val <= 247;
                622 : val <= 247;
                623 : val <= 247;
                624 : val <= 247;
                625 : val <= 247;
                626 : val <= 247;
                627 : val <= 247;
                628 : val <= 247;
                629 : val <= 246;
                630 : val <= 246;
                631 : val <= 246;
                632 : val <= 246;
                633 : val <= 246;
                634 : val <= 246;
                635 : val <= 246;
                636 : val <= 245;
                637 : val <= 245;
                638 : val <= 245;
                639 : val <= 245;
                640 : val <= 245;
                641 : val <= 245;
                642 : val <= 244;
                643 : val <= 244;
                644 : val <= 244;
                645 : val <= 244;
                646 : val <= 244;
                647 : val <= 244;
                648 : val <= 244;
                649 : val <= 243;
                650 : val <= 243;
                651 : val <= 243;
                652 : val <= 243;
                653 : val <= 243;
                654 : val <= 243;
                655 : val <= 242;
                656 : val <= 242;
                657 : val <= 242;
                658 : val <= 242;
                659 : val <= 242;
                660 : val <= 242;
                661 : val <= 241;
                662 : val <= 241;
                663 : val <= 241;
                664 : val <= 241;
                665 : val <= 241;
                666 : val <= 241;
                667 : val <= 240;
                668 : val <= 240;
                669 : val <= 240;
                670 : val <= 240;
                671 : val <= 240;
                672 : val <= 239;
                673 : val <= 239;
                674 : val <= 239;
                675 : val <= 239;
                676 : val <= 239;
                677 : val <= 239;
                678 : val <= 238;
                679 : val <= 238;
                680 : val <= 238;
                681 : val <= 238;
                682 : val <= 238;
                683 : val <= 237;
                684 : val <= 237;
                685 : val <= 237;
                686 : val <= 237;
                687 : val <= 237;
                688 : val <= 236;
                689 : val <= 236;
                690 : val <= 236;
                691 : val <= 236;
                692 : val <= 236;
                693 : val <= 235;
                694 : val <= 235;
                695 : val <= 235;
                696 : val <= 235;
                697 : val <= 235;
                698 : val <= 234;
                699 : val <= 234;
                700 : val <= 234;
                701 : val <= 234;
                702 : val <= 233;
                703 : val <= 233;
                704 : val <= 233;
                705 : val <= 233;
                706 : val <= 233;
                707 : val <= 232;
                708 : val <= 232;
                709 : val <= 232;
                710 : val <= 232;
                711 : val <= 231;
                712 : val <= 231;
                713 : val <= 231;
                714 : val <= 231;
                715 : val <= 231;
                716 : val <= 230;
                717 : val <= 230;
                718 : val <= 230;
                719 : val <= 230;
                720 : val <= 229;
                721 : val <= 229;
                722 : val <= 229;
                723 : val <= 229;
                724 : val <= 228;
                725 : val <= 228;
                726 : val <= 228;
                727 : val <= 228;
                728 : val <= 228;
                729 : val <= 227;
                730 : val <= 227;
                731 : val <= 227;
                732 : val <= 227;
                733 : val <= 226;
                734 : val <= 226;
                735 : val <= 226;
                736 : val <= 226;
                737 : val <= 225;
                738 : val <= 225;
                739 : val <= 225;
                740 : val <= 225;
                741 : val <= 224;
                742 : val <= 224;
                743 : val <= 224;
                744 : val <= 224;
                745 : val <= 223;
                746 : val <= 223;
                747 : val <= 223;
                748 : val <= 223;
                749 : val <= 222;
                750 : val <= 222;
                751 : val <= 222;
                752 : val <= 221;
                753 : val <= 221;
                754 : val <= 221;
                755 : val <= 221;
                756 : val <= 220;
                757 : val <= 220;
                758 : val <= 220;
                759 : val <= 220;
                760 : val <= 219;
                761 : val <= 219;
                762 : val <= 219;
                763 : val <= 219;
                764 : val <= 218;
                765 : val <= 218;
                766 : val <= 218;
                767 : val <= 217;
                768 : val <= 217;
                769 : val <= 217;
                770 : val <= 217;
                771 : val <= 216;
                772 : val <= 216;
                773 : val <= 216;
                774 : val <= 215;
                775 : val <= 215;
                776 : val <= 215;
                777 : val <= 215;
                778 : val <= 214;
                779 : val <= 214;
                780 : val <= 214;
                781 : val <= 213;
                782 : val <= 213;
                783 : val <= 213;
                784 : val <= 213;
                785 : val <= 212;
                786 : val <= 212;
                787 : val <= 212;
                788 : val <= 211;
                789 : val <= 211;
                790 : val <= 211;
                791 : val <= 211;
                792 : val <= 210;
                793 : val <= 210;
                794 : val <= 210;
                795 : val <= 209;
                796 : val <= 209;
                797 : val <= 209;
                798 : val <= 208;
                799 : val <= 208;
                800 : val <= 208;
                801 : val <= 208;
                802 : val <= 207;
                803 : val <= 207;
                804 : val <= 207;
                805 : val <= 206;
                806 : val <= 206;
                807 : val <= 206;
                808 : val <= 205;
                809 : val <= 205;
                810 : val <= 205;
                811 : val <= 205;
                812 : val <= 204;
                813 : val <= 204;
                814 : val <= 204;
                815 : val <= 203;
                816 : val <= 203;
                817 : val <= 203;
                818 : val <= 202;
                819 : val <= 202;
                820 : val <= 202;
                821 : val <= 201;
                822 : val <= 201;
                823 : val <= 201;
                824 : val <= 200;
                825 : val <= 200;
                826 : val <= 200;
                827 : val <= 199;
                828 : val <= 199;
                829 : val <= 199;
                830 : val <= 198;
                831 : val <= 198;
                832 : val <= 198;
                833 : val <= 198;
                834 : val <= 197;
                835 : val <= 197;
                836 : val <= 197;
                837 : val <= 196;
                838 : val <= 196;
                839 : val <= 196;
                840 : val <= 195;
                841 : val <= 195;
                842 : val <= 195;
                843 : val <= 194;
                844 : val <= 194;
                845 : val <= 194;
                846 : val <= 193;
                847 : val <= 193;
                848 : val <= 193;
                849 : val <= 192;
                850 : val <= 192;
                851 : val <= 192;
                852 : val <= 191;
                853 : val <= 191;
                854 : val <= 191;
                855 : val <= 190;
                856 : val <= 190;
                857 : val <= 190;
                858 : val <= 189;
                859 : val <= 189;
                860 : val <= 188;
                861 : val <= 188;
                862 : val <= 188;
                863 : val <= 187;
                864 : val <= 187;
                865 : val <= 187;
                866 : val <= 186;
                867 : val <= 186;
                868 : val <= 186;
                869 : val <= 185;
                870 : val <= 185;
                871 : val <= 185;
                872 : val <= 184;
                873 : val <= 184;
                874 : val <= 184;
                875 : val <= 183;
                876 : val <= 183;
                877 : val <= 183;
                878 : val <= 182;
                879 : val <= 182;
                880 : val <= 182;
                881 : val <= 181;
                882 : val <= 181;
                883 : val <= 180;
                884 : val <= 180;
                885 : val <= 180;
                886 : val <= 179;
                887 : val <= 179;
                888 : val <= 179;
                889 : val <= 178;
                890 : val <= 178;
                891 : val <= 178;
                892 : val <= 177;
                893 : val <= 177;
                894 : val <= 177;
                895 : val <= 176;
                896 : val <= 176;
                897 : val <= 175;
                898 : val <= 175;
                899 : val <= 175;
                900 : val <= 174;
                901 : val <= 174;
                902 : val <= 174;
                903 : val <= 173;
                904 : val <= 173;
                905 : val <= 173;
                906 : val <= 172;
                907 : val <= 172;
                908 : val <= 171;
                909 : val <= 171;
                910 : val <= 171;
                911 : val <= 170;
                912 : val <= 170;
                913 : val <= 170;
                914 : val <= 169;
                915 : val <= 169;
                916 : val <= 168;
                917 : val <= 168;
                918 : val <= 168;
                919 : val <= 167;
                920 : val <= 167;
                921 : val <= 167;
                922 : val <= 166;
                923 : val <= 166;
                924 : val <= 166;
                925 : val <= 165;
                926 : val <= 165;
                927 : val <= 164;
                928 : val <= 164;
                929 : val <= 164;
                930 : val <= 163;
                931 : val <= 163;
                932 : val <= 163;
                933 : val <= 162;
                934 : val <= 162;
                935 : val <= 161;
                936 : val <= 161;
                937 : val <= 161;
                938 : val <= 160;
                939 : val <= 160;
                940 : val <= 159;
                941 : val <= 159;
                942 : val <= 159;
                943 : val <= 158;
                944 : val <= 158;
                945 : val <= 158;
                946 : val <= 157;
                947 : val <= 157;
                948 : val <= 156;
                949 : val <= 156;
                950 : val <= 156;
                951 : val <= 155;
                952 : val <= 155;
                953 : val <= 155;
                954 : val <= 154;
                955 : val <= 154;
                956 : val <= 153;
                957 : val <= 153;
                958 : val <= 153;
                959 : val <= 152;
                960 : val <= 152;
                961 : val <= 151;
                962 : val <= 151;
                963 : val <= 151;
                964 : val <= 150;
                965 : val <= 150;
                966 : val <= 150;
                967 : val <= 149;
                968 : val <= 149;
                969 : val <= 148;
                970 : val <= 148;
                971 : val <= 148;
                972 : val <= 147;
                973 : val <= 147;
                974 : val <= 146;
                975 : val <= 146;
                976 : val <= 146;
                977 : val <= 145;
                978 : val <= 145;
                979 : val <= 145;
                980 : val <= 144;
                981 : val <= 144;
                982 : val <= 143;
                983 : val <= 143;
                984 : val <= 143;
                985 : val <= 142;
                986 : val <= 142;
                987 : val <= 141;
                988 : val <= 141;
                989 : val <= 141;
                990 : val <= 140;
                991 : val <= 140;
                992 : val <= 139;
                993 : val <= 139;
                994 : val <= 139;
                995 : val <= 138;
                996 : val <= 138;
                997 : val <= 138;
                998 : val <= 137;
                999 : val <= 137;
                1000 : val <= 136;
                1001 : val <= 136;
                1002 : val <= 136;
                1003 : val <= 135;
                1004 : val <= 135;
                1005 : val <= 134;
                1006 : val <= 134;
                1007 : val <= 134;
                1008 : val <= 133;
                1009 : val <= 133;
                1010 : val <= 132;
                1011 : val <= 132;
                1012 : val <= 132;
                1013 : val <= 131;
                1014 : val <= 131;
                1015 : val <= 131;
                1016 : val <= 130;
                1017 : val <= 130;
                1018 : val <= 129;
                1019 : val <= 129;
                1020 : val <= 129;
                1021 : val <= 128;
                1022 : val <= 128;
                1023 : val <= 127;
                1024 : val <= 127;
                1025 : val <= 127;
                1026 : val <= 126;
                1027 : val <= 126;
                1028 : val <= 125;
                1029 : val <= 125;
                1030 : val <= 125;
                1031 : val <= 124;
                1032 : val <= 124;
                1033 : val <= 123;
                1034 : val <= 123;
                1035 : val <= 123;
                1036 : val <= 122;
                1037 : val <= 122;
                1038 : val <= 122;
                1039 : val <= 121;
                1040 : val <= 121;
                1041 : val <= 120;
                1042 : val <= 120;
                1043 : val <= 120;
                1044 : val <= 119;
                1045 : val <= 119;
                1046 : val <= 118;
                1047 : val <= 118;
                1048 : val <= 118;
                1049 : val <= 117;
                1050 : val <= 117;
                1051 : val <= 116;
                1052 : val <= 116;
                1053 : val <= 116;
                1054 : val <= 115;
                1055 : val <= 115;
                1056 : val <= 115;
                1057 : val <= 114;
                1058 : val <= 114;
                1059 : val <= 113;
                1060 : val <= 113;
                1061 : val <= 113;
                1062 : val <= 112;
                1063 : val <= 112;
                1064 : val <= 111;
                1065 : val <= 111;
                1066 : val <= 111;
                1067 : val <= 110;
                1068 : val <= 110;
                1069 : val <= 109;
                1070 : val <= 109;
                1071 : val <= 109;
                1072 : val <= 108;
                1073 : val <= 108;
                1074 : val <= 108;
                1075 : val <= 107;
                1076 : val <= 107;
                1077 : val <= 106;
                1078 : val <= 106;
                1079 : val <= 106;
                1080 : val <= 105;
                1081 : val <= 105;
                1082 : val <= 104;
                1083 : val <= 104;
                1084 : val <= 104;
                1085 : val <= 103;
                1086 : val <= 103;
                1087 : val <= 103;
                1088 : val <= 102;
                1089 : val <= 102;
                1090 : val <= 101;
                1091 : val <= 101;
                1092 : val <= 101;
                1093 : val <= 100;
                1094 : val <= 100;
                1095 : val <= 99;
                1096 : val <= 99;
                1097 : val <= 99;
                1098 : val <= 98;
                1099 : val <= 98;
                1100 : val <= 98;
                1101 : val <= 97;
                1102 : val <= 97;
                1103 : val <= 96;
                1104 : val <= 96;
                1105 : val <= 96;
                1106 : val <= 95;
                1107 : val <= 95;
                1108 : val <= 95;
                1109 : val <= 94;
                1110 : val <= 94;
                1111 : val <= 93;
                1112 : val <= 93;
                1113 : val <= 93;
                1114 : val <= 92;
                1115 : val <= 92;
                1116 : val <= 91;
                1117 : val <= 91;
                1118 : val <= 91;
                1119 : val <= 90;
                1120 : val <= 90;
                1121 : val <= 90;
                1122 : val <= 89;
                1123 : val <= 89;
                1124 : val <= 88;
                1125 : val <= 88;
                1126 : val <= 88;
                1127 : val <= 87;
                1128 : val <= 87;
                1129 : val <= 87;
                1130 : val <= 86;
                1131 : val <= 86;
                1132 : val <= 86;
                1133 : val <= 85;
                1134 : val <= 85;
                1135 : val <= 84;
                1136 : val <= 84;
                1137 : val <= 84;
                1138 : val <= 83;
                1139 : val <= 83;
                1140 : val <= 83;
                1141 : val <= 82;
                1142 : val <= 82;
                1143 : val <= 81;
                1144 : val <= 81;
                1145 : val <= 81;
                1146 : val <= 80;
                1147 : val <= 80;
                1148 : val <= 80;
                1149 : val <= 79;
                1150 : val <= 79;
                1151 : val <= 79;
                1152 : val <= 78;
                1153 : val <= 78;
                1154 : val <= 77;
                1155 : val <= 77;
                1156 : val <= 77;
                1157 : val <= 76;
                1158 : val <= 76;
                1159 : val <= 76;
                1160 : val <= 75;
                1161 : val <= 75;
                1162 : val <= 75;
                1163 : val <= 74;
                1164 : val <= 74;
                1165 : val <= 74;
                1166 : val <= 73;
                1167 : val <= 73;
                1168 : val <= 72;
                1169 : val <= 72;
                1170 : val <= 72;
                1171 : val <= 71;
                1172 : val <= 71;
                1173 : val <= 71;
                1174 : val <= 70;
                1175 : val <= 70;
                1176 : val <= 70;
                1177 : val <= 69;
                1178 : val <= 69;
                1179 : val <= 69;
                1180 : val <= 68;
                1181 : val <= 68;
                1182 : val <= 68;
                1183 : val <= 67;
                1184 : val <= 67;
                1185 : val <= 67;
                1186 : val <= 66;
                1187 : val <= 66;
                1188 : val <= 66;
                1189 : val <= 65;
                1190 : val <= 65;
                1191 : val <= 64;
                1192 : val <= 64;
                1193 : val <= 64;
                1194 : val <= 63;
                1195 : val <= 63;
                1196 : val <= 63;
                1197 : val <= 62;
                1198 : val <= 62;
                1199 : val <= 62;
                1200 : val <= 61;
                1201 : val <= 61;
                1202 : val <= 61;
                1203 : val <= 60;
                1204 : val <= 60;
                1205 : val <= 60;
                1206 : val <= 59;
                1207 : val <= 59;
                1208 : val <= 59;
                1209 : val <= 58;
                1210 : val <= 58;
                1211 : val <= 58;
                1212 : val <= 57;
                1213 : val <= 57;
                1214 : val <= 57;
                1215 : val <= 56;
                1216 : val <= 56;
                1217 : val <= 56;
                1218 : val <= 56;
                1219 : val <= 55;
                1220 : val <= 55;
                1221 : val <= 55;
                1222 : val <= 54;
                1223 : val <= 54;
                1224 : val <= 54;
                1225 : val <= 53;
                1226 : val <= 53;
                1227 : val <= 53;
                1228 : val <= 52;
                1229 : val <= 52;
                1230 : val <= 52;
                1231 : val <= 51;
                1232 : val <= 51;
                1233 : val <= 51;
                1234 : val <= 50;
                1235 : val <= 50;
                1236 : val <= 50;
                1237 : val <= 49;
                1238 : val <= 49;
                1239 : val <= 49;
                1240 : val <= 49;
                1241 : val <= 48;
                1242 : val <= 48;
                1243 : val <= 48;
                1244 : val <= 47;
                1245 : val <= 47;
                1246 : val <= 47;
                1247 : val <= 46;
                1248 : val <= 46;
                1249 : val <= 46;
                1250 : val <= 46;
                1251 : val <= 45;
                1252 : val <= 45;
                1253 : val <= 45;
                1254 : val <= 44;
                1255 : val <= 44;
                1256 : val <= 44;
                1257 : val <= 43;
                1258 : val <= 43;
                1259 : val <= 43;
                1260 : val <= 43;
                1261 : val <= 42;
                1262 : val <= 42;
                1263 : val <= 42;
                1264 : val <= 41;
                1265 : val <= 41;
                1266 : val <= 41;
                1267 : val <= 41;
                1268 : val <= 40;
                1269 : val <= 40;
                1270 : val <= 40;
                1271 : val <= 39;
                1272 : val <= 39;
                1273 : val <= 39;
                1274 : val <= 39;
                1275 : val <= 38;
                1276 : val <= 38;
                1277 : val <= 38;
                1278 : val <= 37;
                1279 : val <= 37;
                1280 : val <= 37;
                1281 : val <= 37;
                1282 : val <= 36;
                1283 : val <= 36;
                1284 : val <= 36;
                1285 : val <= 35;
                1286 : val <= 35;
                1287 : val <= 35;
                1288 : val <= 35;
                1289 : val <= 34;
                1290 : val <= 34;
                1291 : val <= 34;
                1292 : val <= 34;
                1293 : val <= 33;
                1294 : val <= 33;
                1295 : val <= 33;
                1296 : val <= 33;
                1297 : val <= 32;
                1298 : val <= 32;
                1299 : val <= 32;
                1300 : val <= 31;
                1301 : val <= 31;
                1302 : val <= 31;
                1303 : val <= 31;
                1304 : val <= 30;
                1305 : val <= 30;
                1306 : val <= 30;
                1307 : val <= 30;
                1308 : val <= 29;
                1309 : val <= 29;
                1310 : val <= 29;
                1311 : val <= 29;
                1312 : val <= 28;
                1313 : val <= 28;
                1314 : val <= 28;
                1315 : val <= 28;
                1316 : val <= 27;
                1317 : val <= 27;
                1318 : val <= 27;
                1319 : val <= 27;
                1320 : val <= 26;
                1321 : val <= 26;
                1322 : val <= 26;
                1323 : val <= 26;
                1324 : val <= 26;
                1325 : val <= 25;
                1326 : val <= 25;
                1327 : val <= 25;
                1328 : val <= 25;
                1329 : val <= 24;
                1330 : val <= 24;
                1331 : val <= 24;
                1332 : val <= 24;
                1333 : val <= 23;
                1334 : val <= 23;
                1335 : val <= 23;
                1336 : val <= 23;
                1337 : val <= 23;
                1338 : val <= 22;
                1339 : val <= 22;
                1340 : val <= 22;
                1341 : val <= 22;
                1342 : val <= 21;
                1343 : val <= 21;
                1344 : val <= 21;
                1345 : val <= 21;
                1346 : val <= 21;
                1347 : val <= 20;
                1348 : val <= 20;
                1349 : val <= 20;
                1350 : val <= 20;
                1351 : val <= 19;
                1352 : val <= 19;
                1353 : val <= 19;
                1354 : val <= 19;
                1355 : val <= 19;
                1356 : val <= 18;
                1357 : val <= 18;
                1358 : val <= 18;
                1359 : val <= 18;
                1360 : val <= 18;
                1361 : val <= 17;
                1362 : val <= 17;
                1363 : val <= 17;
                1364 : val <= 17;
                1365 : val <= 17;
                1366 : val <= 16;
                1367 : val <= 16;
                1368 : val <= 16;
                1369 : val <= 16;
                1370 : val <= 16;
                1371 : val <= 15;
                1372 : val <= 15;
                1373 : val <= 15;
                1374 : val <= 15;
                1375 : val <= 15;
                1376 : val <= 15;
                1377 : val <= 14;
                1378 : val <= 14;
                1379 : val <= 14;
                1380 : val <= 14;
                1381 : val <= 14;
                1382 : val <= 13;
                1383 : val <= 13;
                1384 : val <= 13;
                1385 : val <= 13;
                1386 : val <= 13;
                1387 : val <= 13;
                1388 : val <= 12;
                1389 : val <= 12;
                1390 : val <= 12;
                1391 : val <= 12;
                1392 : val <= 12;
                1393 : val <= 12;
                1394 : val <= 11;
                1395 : val <= 11;
                1396 : val <= 11;
                1397 : val <= 11;
                1398 : val <= 11;
                1399 : val <= 11;
                1400 : val <= 10;
                1401 : val <= 10;
                1402 : val <= 10;
                1403 : val <= 10;
                1404 : val <= 10;
                1405 : val <= 10;
                1406 : val <= 10;
                1407 : val <= 9;
                1408 : val <= 9;
                1409 : val <= 9;
                1410 : val <= 9;
                1411 : val <= 9;
                1412 : val <= 9;
                1413 : val <= 8;
                1414 : val <= 8;
                1415 : val <= 8;
                1416 : val <= 8;
                1417 : val <= 8;
                1418 : val <= 8;
                1419 : val <= 8;
                1420 : val <= 7;
                1421 : val <= 7;
                1422 : val <= 7;
                1423 : val <= 7;
                1424 : val <= 7;
                1425 : val <= 7;
                1426 : val <= 7;
                1427 : val <= 7;
                1428 : val <= 6;
                1429 : val <= 6;
                1430 : val <= 6;
                1431 : val <= 6;
                1432 : val <= 6;
                1433 : val <= 6;
                1434 : val <= 6;
                1435 : val <= 6;
                1436 : val <= 5;
                1437 : val <= 5;
                1438 : val <= 5;
                1439 : val <= 5;
                1440 : val <= 5;
                1441 : val <= 5;
                1442 : val <= 5;
                1443 : val <= 5;
                1444 : val <= 5;
                1445 : val <= 4;
                1446 : val <= 4;
                1447 : val <= 4;
                1448 : val <= 4;
                1449 : val <= 4;
                1450 : val <= 4;
                1451 : val <= 4;
                1452 : val <= 4;
                1453 : val <= 4;
                1454 : val <= 4;
                1455 : val <= 3;
                1456 : val <= 3;
                1457 : val <= 3;
                1458 : val <= 3;
                1459 : val <= 3;
                1460 : val <= 3;
                1461 : val <= 3;
                1462 : val <= 3;
                1463 : val <= 3;
                1464 : val <= 3;
                1465 : val <= 3;
                1466 : val <= 2;
                1467 : val <= 2;
                1468 : val <= 2;
                1469 : val <= 2;
                1470 : val <= 2;
                1471 : val <= 2;
                1472 : val <= 2;
                1473 : val <= 2;
                1474 : val <= 2;
                1475 : val <= 2;
                1476 : val <= 2;
                1477 : val <= 2;
                1478 : val <= 2;
                1479 : val <= 1;
                1480 : val <= 1;
                1481 : val <= 1;
                1482 : val <= 1;
                1483 : val <= 1;
                1484 : val <= 1;
                1485 : val <= 1;
                1486 : val <= 1;
                1487 : val <= 1;
                1488 : val <= 1;
                1489 : val <= 1;
                1490 : val <= 1;
                1491 : val <= 1;
                1492 : val <= 1;
                1493 : val <= 1;
                1494 : val <= 1;
                1495 : val <= 1;
                1496 : val <= 0;
                1497 : val <= 0;
                1498 : val <= 0;
                1499 : val <= 0;
                1500 : val <= 0;
                1501 : val <= 0;
                1502 : val <= 0;
                1503 : val <= 0;
                1504 : val <= 0;
                1505 : val <= 0;
                1506 : val <= 0;
                1507 : val <= 0;
                1508 : val <= 0;
                1509 : val <= 0;
                1510 : val <= 0;
                1511 : val <= 0;
                1512 : val <= 0;
                1513 : val <= 0;
                1514 : val <= 0;
                1515 : val <= 0;
                1516 : val <= 0;
                1517 : val <= 0;
                1518 : val <= 0;
                1519 : val <= 0;
                1520 : val <= 0;
                1521 : val <= 0;
                1522 : val <= 0;
                1523 : val <= 0;
                1524 : val <= 0;
                1525 : val <= 0;
                1526 : val <= 0;
                1527 : val <= 0;
                1528 : val <= 0;
                1529 : val <= 0;
                1530 : val <= 0;
                1531 : val <= 0;
                1532 : val <= 0;
                1533 : val <= 0;
                1534 : val <= 0;
                1535 : val <= 0;
                1536 : val <= -1;
                1537 : val <= 0;
                1538 : val <= 0;
                1539 : val <= 0;
                1540 : val <= 0;
                1541 : val <= 0;
                1542 : val <= 0;
                1543 : val <= 0;
                1544 : val <= 0;
                1545 : val <= 0;
                1546 : val <= 0;
                1547 : val <= 0;
                1548 : val <= 0;
                1549 : val <= 0;
                1550 : val <= 0;
                1551 : val <= 0;
                1552 : val <= 0;
                1553 : val <= 0;
                1554 : val <= 0;
                1555 : val <= 0;
                1556 : val <= 0;
                1557 : val <= 0;
                1558 : val <= 0;
                1559 : val <= 0;
                1560 : val <= 0;
                1561 : val <= 0;
                1562 : val <= 0;
                1563 : val <= 0;
                1564 : val <= 0;
                1565 : val <= 0;
                1566 : val <= 0;
                1567 : val <= 0;
                1568 : val <= 0;
                1569 : val <= 0;
                1570 : val <= 0;
                1571 : val <= 0;
                1572 : val <= 0;
                1573 : val <= 0;
                1574 : val <= 0;
                1575 : val <= 0;
                1576 : val <= 0;
                1577 : val <= 1;
                1578 : val <= 1;
                1579 : val <= 1;
                1580 : val <= 1;
                1581 : val <= 1;
                1582 : val <= 1;
                1583 : val <= 1;
                1584 : val <= 1;
                1585 : val <= 1;
                1586 : val <= 1;
                1587 : val <= 1;
                1588 : val <= 1;
                1589 : val <= 1;
                1590 : val <= 1;
                1591 : val <= 1;
                1592 : val <= 1;
                1593 : val <= 1;
                1594 : val <= 2;
                1595 : val <= 2;
                1596 : val <= 2;
                1597 : val <= 2;
                1598 : val <= 2;
                1599 : val <= 2;
                1600 : val <= 2;
                1601 : val <= 2;
                1602 : val <= 2;
                1603 : val <= 2;
                1604 : val <= 2;
                1605 : val <= 2;
                1606 : val <= 2;
                1607 : val <= 3;
                1608 : val <= 3;
                1609 : val <= 3;
                1610 : val <= 3;
                1611 : val <= 3;
                1612 : val <= 3;
                1613 : val <= 3;
                1614 : val <= 3;
                1615 : val <= 3;
                1616 : val <= 3;
                1617 : val <= 3;
                1618 : val <= 4;
                1619 : val <= 4;
                1620 : val <= 4;
                1621 : val <= 4;
                1622 : val <= 4;
                1623 : val <= 4;
                1624 : val <= 4;
                1625 : val <= 4;
                1626 : val <= 4;
                1627 : val <= 4;
                1628 : val <= 5;
                1629 : val <= 5;
                1630 : val <= 5;
                1631 : val <= 5;
                1632 : val <= 5;
                1633 : val <= 5;
                1634 : val <= 5;
                1635 : val <= 5;
                1636 : val <= 5;
                1637 : val <= 6;
                1638 : val <= 6;
                1639 : val <= 6;
                1640 : val <= 6;
                1641 : val <= 6;
                1642 : val <= 6;
                1643 : val <= 6;
                1644 : val <= 6;
                1645 : val <= 7;
                1646 : val <= 7;
                1647 : val <= 7;
                1648 : val <= 7;
                1649 : val <= 7;
                1650 : val <= 7;
                1651 : val <= 7;
                1652 : val <= 7;
                1653 : val <= 8;
                1654 : val <= 8;
                1655 : val <= 8;
                1656 : val <= 8;
                1657 : val <= 8;
                1658 : val <= 8;
                1659 : val <= 8;
                1660 : val <= 9;
                1661 : val <= 9;
                1662 : val <= 9;
                1663 : val <= 9;
                1664 : val <= 9;
                1665 : val <= 9;
                1666 : val <= 10;
                1667 : val <= 10;
                1668 : val <= 10;
                1669 : val <= 10;
                1670 : val <= 10;
                1671 : val <= 10;
                1672 : val <= 10;
                1673 : val <= 11;
                1674 : val <= 11;
                1675 : val <= 11;
                1676 : val <= 11;
                1677 : val <= 11;
                1678 : val <= 11;
                1679 : val <= 12;
                1680 : val <= 12;
                1681 : val <= 12;
                1682 : val <= 12;
                1683 : val <= 12;
                1684 : val <= 12;
                1685 : val <= 13;
                1686 : val <= 13;
                1687 : val <= 13;
                1688 : val <= 13;
                1689 : val <= 13;
                1690 : val <= 13;
                1691 : val <= 14;
                1692 : val <= 14;
                1693 : val <= 14;
                1694 : val <= 14;
                1695 : val <= 14;
                1696 : val <= 15;
                1697 : val <= 15;
                1698 : val <= 15;
                1699 : val <= 15;
                1700 : val <= 15;
                1701 : val <= 15;
                1702 : val <= 16;
                1703 : val <= 16;
                1704 : val <= 16;
                1705 : val <= 16;
                1706 : val <= 16;
                1707 : val <= 17;
                1708 : val <= 17;
                1709 : val <= 17;
                1710 : val <= 17;
                1711 : val <= 17;
                1712 : val <= 18;
                1713 : val <= 18;
                1714 : val <= 18;
                1715 : val <= 18;
                1716 : val <= 18;
                1717 : val <= 19;
                1718 : val <= 19;
                1719 : val <= 19;
                1720 : val <= 19;
                1721 : val <= 19;
                1722 : val <= 20;
                1723 : val <= 20;
                1724 : val <= 20;
                1725 : val <= 20;
                1726 : val <= 21;
                1727 : val <= 21;
                1728 : val <= 21;
                1729 : val <= 21;
                1730 : val <= 21;
                1731 : val <= 22;
                1732 : val <= 22;
                1733 : val <= 22;
                1734 : val <= 22;
                1735 : val <= 23;
                1736 : val <= 23;
                1737 : val <= 23;
                1738 : val <= 23;
                1739 : val <= 23;
                1740 : val <= 24;
                1741 : val <= 24;
                1742 : val <= 24;
                1743 : val <= 24;
                1744 : val <= 25;
                1745 : val <= 25;
                1746 : val <= 25;
                1747 : val <= 25;
                1748 : val <= 26;
                1749 : val <= 26;
                1750 : val <= 26;
                1751 : val <= 26;
                1752 : val <= 26;
                1753 : val <= 27;
                1754 : val <= 27;
                1755 : val <= 27;
                1756 : val <= 27;
                1757 : val <= 28;
                1758 : val <= 28;
                1759 : val <= 28;
                1760 : val <= 28;
                1761 : val <= 29;
                1762 : val <= 29;
                1763 : val <= 29;
                1764 : val <= 29;
                1765 : val <= 30;
                1766 : val <= 30;
                1767 : val <= 30;
                1768 : val <= 30;
                1769 : val <= 31;
                1770 : val <= 31;
                1771 : val <= 31;
                1772 : val <= 31;
                1773 : val <= 32;
                1774 : val <= 32;
                1775 : val <= 32;
                1776 : val <= 33;
                1777 : val <= 33;
                1778 : val <= 33;
                1779 : val <= 33;
                1780 : val <= 34;
                1781 : val <= 34;
                1782 : val <= 34;
                1783 : val <= 34;
                1784 : val <= 35;
                1785 : val <= 35;
                1786 : val <= 35;
                1787 : val <= 35;
                1788 : val <= 36;
                1789 : val <= 36;
                1790 : val <= 36;
                1791 : val <= 37;
                1792 : val <= 37;
                1793 : val <= 37;
                1794 : val <= 37;
                1795 : val <= 38;
                1796 : val <= 38;
                1797 : val <= 38;
                1798 : val <= 39;
                1799 : val <= 39;
                1800 : val <= 39;
                1801 : val <= 39;
                1802 : val <= 40;
                1803 : val <= 40;
                1804 : val <= 40;
                1805 : val <= 41;
                1806 : val <= 41;
                1807 : val <= 41;
                1808 : val <= 41;
                1809 : val <= 42;
                1810 : val <= 42;
                1811 : val <= 42;
                1812 : val <= 43;
                1813 : val <= 43;
                1814 : val <= 43;
                1815 : val <= 43;
                1816 : val <= 44;
                1817 : val <= 44;
                1818 : val <= 44;
                1819 : val <= 45;
                1820 : val <= 45;
                1821 : val <= 45;
                1822 : val <= 46;
                1823 : val <= 46;
                1824 : val <= 46;
                1825 : val <= 46;
                1826 : val <= 47;
                1827 : val <= 47;
                1828 : val <= 47;
                1829 : val <= 48;
                1830 : val <= 48;
                1831 : val <= 48;
                1832 : val <= 49;
                1833 : val <= 49;
                1834 : val <= 49;
                1835 : val <= 49;
                1836 : val <= 50;
                1837 : val <= 50;
                1838 : val <= 50;
                1839 : val <= 51;
                1840 : val <= 51;
                1841 : val <= 51;
                1842 : val <= 52;
                1843 : val <= 52;
                1844 : val <= 52;
                1845 : val <= 53;
                1846 : val <= 53;
                1847 : val <= 53;
                1848 : val <= 54;
                1849 : val <= 54;
                1850 : val <= 54;
                1851 : val <= 55;
                1852 : val <= 55;
                1853 : val <= 55;
                1854 : val <= 56;
                1855 : val <= 56;
                1856 : val <= 56;
                1857 : val <= 56;
                1858 : val <= 57;
                1859 : val <= 57;
                1860 : val <= 57;
                1861 : val <= 58;
                1862 : val <= 58;
                1863 : val <= 58;
                1864 : val <= 59;
                1865 : val <= 59;
                1866 : val <= 59;
                1867 : val <= 60;
                1868 : val <= 60;
                1869 : val <= 60;
                1870 : val <= 61;
                1871 : val <= 61;
                1872 : val <= 61;
                1873 : val <= 62;
                1874 : val <= 62;
                1875 : val <= 62;
                1876 : val <= 63;
                1877 : val <= 63;
                1878 : val <= 63;
                1879 : val <= 64;
                1880 : val <= 64;
                1881 : val <= 64;
                1882 : val <= 65;
                1883 : val <= 65;
                1884 : val <= 66;
                1885 : val <= 66;
                1886 : val <= 66;
                1887 : val <= 67;
                1888 : val <= 67;
                1889 : val <= 67;
                1890 : val <= 68;
                1891 : val <= 68;
                1892 : val <= 68;
                1893 : val <= 69;
                1894 : val <= 69;
                1895 : val <= 69;
                1896 : val <= 70;
                1897 : val <= 70;
                1898 : val <= 70;
                1899 : val <= 71;
                1900 : val <= 71;
                1901 : val <= 71;
                1902 : val <= 72;
                1903 : val <= 72;
                1904 : val <= 72;
                1905 : val <= 73;
                1906 : val <= 73;
                1907 : val <= 74;
                1908 : val <= 74;
                1909 : val <= 74;
                1910 : val <= 75;
                1911 : val <= 75;
                1912 : val <= 75;
                1913 : val <= 76;
                1914 : val <= 76;
                1915 : val <= 76;
                1916 : val <= 77;
                1917 : val <= 77;
                1918 : val <= 77;
                1919 : val <= 78;
                1920 : val <= 78;
                1921 : val <= 79;
                1922 : val <= 79;
                1923 : val <= 79;
                1924 : val <= 80;
                1925 : val <= 80;
                1926 : val <= 80;
                1927 : val <= 81;
                1928 : val <= 81;
                1929 : val <= 81;
                1930 : val <= 82;
                1931 : val <= 82;
                1932 : val <= 83;
                1933 : val <= 83;
                1934 : val <= 83;
                1935 : val <= 84;
                1936 : val <= 84;
                1937 : val <= 84;
                1938 : val <= 85;
                1939 : val <= 85;
                1940 : val <= 86;
                1941 : val <= 86;
                1942 : val <= 86;
                1943 : val <= 87;
                1944 : val <= 87;
                1945 : val <= 87;
                1946 : val <= 88;
                1947 : val <= 88;
                1948 : val <= 88;
                1949 : val <= 89;
                1950 : val <= 89;
                1951 : val <= 90;
                1952 : val <= 90;
                1953 : val <= 90;
                1954 : val <= 91;
                1955 : val <= 91;
                1956 : val <= 91;
                1957 : val <= 92;
                1958 : val <= 92;
                1959 : val <= 93;
                1960 : val <= 93;
                1961 : val <= 93;
                1962 : val <= 94;
                1963 : val <= 94;
                1964 : val <= 95;
                1965 : val <= 95;
                1966 : val <= 95;
                1967 : val <= 96;
                1968 : val <= 96;
                1969 : val <= 96;
                1970 : val <= 97;
                1971 : val <= 97;
                1972 : val <= 98;
                1973 : val <= 98;
                1974 : val <= 98;
                1975 : val <= 99;
                1976 : val <= 99;
                1977 : val <= 99;
                1978 : val <= 100;
                1979 : val <= 100;
                1980 : val <= 101;
                1981 : val <= 101;
                1982 : val <= 101;
                1983 : val <= 102;
                1984 : val <= 102;
                1985 : val <= 103;
                1986 : val <= 103;
                1987 : val <= 103;
                1988 : val <= 104;
                1989 : val <= 104;
                1990 : val <= 104;
                1991 : val <= 105;
                1992 : val <= 105;
                1993 : val <= 106;
                1994 : val <= 106;
                1995 : val <= 106;
                1996 : val <= 107;
                1997 : val <= 107;
                1998 : val <= 108;
                1999 : val <= 108;
                2000 : val <= 108;
                2001 : val <= 109;
                2002 : val <= 109;
                2003 : val <= 109;
                2004 : val <= 110;
                2005 : val <= 110;
                2006 : val <= 111;
                2007 : val <= 111;
                2008 : val <= 111;
                2009 : val <= 112;
                2010 : val <= 112;
                2011 : val <= 113;
                2012 : val <= 113;
                2013 : val <= 113;
                2014 : val <= 114;
                2015 : val <= 114;
                2016 : val <= 115;
                2017 : val <= 115;
                2018 : val <= 115;
                2019 : val <= 116;
                2020 : val <= 116;
                2021 : val <= 116;
                2022 : val <= 117;
                2023 : val <= 117;
                2024 : val <= 118;
                2025 : val <= 118;
                2026 : val <= 118;
                2027 : val <= 119;
                2028 : val <= 119;
                2029 : val <= 120;
                2030 : val <= 120;
                2031 : val <= 120;
                2032 : val <= 121;
                2033 : val <= 121;
                2034 : val <= 122;
                2035 : val <= 122;
                2036 : val <= 122;
                2037 : val <= 123;
                2038 : val <= 123;
                2039 : val <= 123;
                2040 : val <= 124;
                2041 : val <= 124;
                2042 : val <= 125;
                2043 : val <= 125;
                2044 : val <= 125;
                2045 : val <= 126;
                2046 : val <= 126;
                2047 : val <= 127;
        endcase

endmodule

