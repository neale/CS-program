module ROM(

	input logic [7:0] buttons,
	input         		encoder0,
	input         		encoder1,
	input         		clk,
	input  wire   		reset,
	input logic       d_out,
	output logic      d_in,
	output 				_sclk,
	output [6:0]  		segments,
	output            dp,
	output [2:0]  		select,
	output 		  		display_clk, //5000Hz
	output        		pwm
	

);
// ADC vars
logic cs_n = 1;
logic [11:0] adc_rom_out;
logic [11:0] d_out_buffer;
logic [3:0]  count_posedge;
logic [3:0]  count_negedge;
logic encoder_a;
logic encoder_b;
logic button0;
logic button1;

// 10K clock
frame_rate frame_rate0(
  .inclk0 ( clk ),
  .c1     ( display_clk ),
  .locked ( lock_display )
);

ADC ADC0 (
	.address ( d_out_buffer ),
	.clock ( _sclk ),
	.q ( adc_rom_out )
);


sclk	sclk_0 (
	.inclk0 ( clk ),
	.c0 ( _sclk )
);

// debounce both of the encoder inputs
debounce encodera(

	.clk       (clk),
	.A		     (encoder0),
	.triggered (encoder_a)
);

debounce encoderb(

	.clk       (clk),
	.A		     (encoder1),
	.triggered (encoder_b)
);

// The adc is free running (may change) at a 2MHZ clk. It has an operating sclk range of 0.8 to 3.2 MHz
// There is a 16 bit data loop that is captured one bit at a time, at the falling edge of sclk
// CS is lowered on the first falling edge, and din is provided one bit at a time at the negedge of sclk
// sclk is raised on the last rising edge of a frame
always @(negedge _sclk)
	begin
   casez(count_negedge)
		
			0 : cs_n = 0;
			2 : d_in = 0;
			3 : d_in = 0;
			4 : d_in = 0;
			default : d_in = 0;
	endcase
	count_negedge++;	
	end
	
always @(posedge _sclk)
	begin
		casez(count_posedge)
			
			4 : d_out_buffer[11] = d_out;
			5 : d_out_buffer[10] = d_out;
			6 : d_out_buffer[9] = d_out;
			7 : d_out_buffer[8] = d_out;
			8 : d_out_buffer[7] = d_out;
			9 : d_out_buffer[6] = d_out;
			10 : d_out_buffer[5] = d_out;
			11 : d_out_buffer[4] = d_out;
			12 : d_out_buffer[3] = d_out;
			13 : d_out_buffer[2] = d_out;
			14 : d_out_buffer[1] = d_out;
			15 : 
				begin
					cs_n = 1;
					d_out_buffer[0] = d_out;
				end
			default : d_out_buffer = 0;
		endcase
		count_posedge++;	
			
	end

// ***************************************************************************//
//										 Routine Logic
// **************************************************************************//
logic [3:0]   digit  = 0;  // initial digit to display

// seven seg decoder
always_comb
	begin
		unique casez (digit)       //abcdefg
										 
			1 : segments = 7'b1111001; 
			2 : segments = 7'b0100100; 
			3 : segments = 7'b0110000; 
			4 : segments = 7'b0011001; 
			5 : segments = 7'b0010010; 
			6 : segments = 7'b0000010; 
			7 : segments = 7'b1111000; 
			8 : segments = 7'b0000000; 
			9 : segments = 7'b0010000; 
			0 : segments = 7'b1000000; 	
			10 : segments = 7'b1111111;
		endcase
	end

// quad encoder logic, Roger';s flip flop idea found on FPGAs are fun
// Takes the known last states of the encoders and debounces them
// Xors a 4 bit register with itself to check for a turn
logic [2:0] encoder0_last;
logic [2:0] encoder1_last;

// sync encoders to the clock
// append encoder states to last states to debounce
// then xor to get final state
always @(posedge clk)
	begin 
		encoder0_last <= {encoder0_last[1:0], encoder_a};
	end
always @(posedge clk)
	begin
		encoder1_last <= {encoder1_last[1:0], encoder_b};
	end
	
wire encoder_turning = encoder0_last[1] ^ encoder0_last[2] ^ encoder1_last[1] ^ encoder1_last[2];
wire encoder_dir   = encoder0_last[1] ^ encoder1_last[2];

// check encoder states, if forward, count up, if backward, count down. 
// count var is 10 bits wide to allow 999 digits
logic [13:0] cnt = 1000;
always  @(posedge clk)
	begin
		if (encoder_turning)
			begin
				if(encoder_dir) 
					cnt<=cnt+1; 
				else 
					cnt<=cnt-1;
				if (cnt > 9999)
					cnt <= cnt - 9999;
			end
		else
			cnt <= cnt;
	end
	
logic [2:0]  select_state = 3'b001;

// state machine for cycling through select_states
// current select bit becomes new select bits
always_ff @ (posedge display_clk)

	begin
		unique casez (select_state)
			3'b001  : select_state = 3'b010; 
			3'b010  : select_state = 3'b100;
			3'b100  : select_state = 3'b111;
			3'b111  : select_state = 3'b001;
		endcase
	end
	
//state machine for cycling through digits
logic [3:0] ones = 0;
logic [3:0] tenth = 0;
logic [3:0] hundredth = 0;
integer  i;
// block takes the current countand creates the digit to push out the decoder
// to do this, we're going to take the 10 bit count value and do some math

//BCD algorithm: double dabble
//or shift and add 3 algorithm

always @ (adc_rom_out)
	begin
        hundredth = 4'd0;
        tenth = 4'd0;
        ones = 4'd0;
		for  (i = 11; i >= 0; i = i-1)
			begin
			  // if the value contained is over 5, add three
			  // so that the shift guarantees the carryover to the next "number"
          if (hundredth >= 5)
               hundredth = hundredth + 3;
			 else
				   hundredth = hundredth;
          if (tenth >= 5)
               tenth = tenth + 3;
			 else
					tenth = tenth;
          if (ones >= 5)
				ones = ones + 3;
			 else
				ones = ones;
			 

          hundredth = hundredth << 1;
          hundredth[0] = tenth[3];
          tenth = tenth << 1;
          tenth[0] = ones[3];
          ones = ones << 1;
          ones[0] = adc_rom_out[i];
				
			end
	end
	
always_comb
	begin
		casez (select)
			3'b011 : dp = 0;
			default: dp = 1;
		endcase
	end
	
always_comb
	begin
	unique casez(select)
		3'b100 : digit = ones; 
		3'b011 : digit = 10;	//always DP on		
		3'b001 : digit = tenth;
		3'b000 : digit = hundredth;
	endcase
	
	end
endmodule
